module Ram (
    input    [6:0]    addr,
    inout    [31:0]    data,
    input              wre,
	 input				  flag,	//memoria de dados/memoria de instrucoes
	 input 				  reset
);

    reg     [31:0]  memory    [0:127];
	 reg     [7:0] i;
	 reg     [7:0] j;

    assign data[31:0] = wre ? memory[addr] : 32'hZZZZ_ZZZZ;

    always @(wre or addr or data or reset) begin
        if (!wre)
            memory[addr] = data[31:0];
				
			if(!reset) begin
				if(flag)begin			
				
					for (i = 8'b0000_1111; i < 128; i = i + 8'b00000001) begin
						memory[i] <= 32'h0000_0000;
					end
					
					memory[0] <= 32'b00100000000000000000000000000001;
					memory[1] <= 32'b00100000001000010000000000000010;// SW,$8,0($0)
					memory[2] <= 32'b00000000000000010001000000100000;
					memory[3] <= 32'b10101100000000100000000000000000;
					memory[4] <= 32'b00000000000000000000000000000000;
					memory[5] <= 32'b00000000000000000000000000000000;
					memory[6] <= 32'b00000000000000000000000000000000;
					memory[7] <= 32'b00000000000000000000000000000000;
					memory[8] <= 32'b00000000000000000000000000000000;
					memory[9] <= 32'b00000000000000000000000000000000;
					/*memory[0] <= 32'b00100001001010010000000000000001;
					memory[1] <= 32'b00100001010010100000000000000010;
					memory[2] <= 32'b00000000000000000000000000000000;
					memory[3] <= 32'b00000001001010100101100000100000;
					memory[4] <= 32'b00000000000000000000000000000000;
					memory[5] <= 32'b00000000000000000000000000000000;
					memory[6] <= 32'b00000001011010100110000000100000;
					memory[9] <= 32'b00000000000000000000000000000000;*/
					memory[10] <= 32'b10001100000000000000000000000000;
				 /*memory[0] <= 32'b001000_00001_00001_0000000000000001;
					memory[1] <= 32'b001000_00010_00010_0000000000000001;
					memory[2] <= 32'b001000_00011_00011_0000000000000100;
					memory[3] <= 32'b000000_00011_00010_00100_00000_011000;
					memory[4] <= 32'b00000000000000000000000000000000;
					memory[5] <= 32'b00000000000000000000000000000000;
					memory[6] <= 32'b00000000000000000000000000000000;
					memory[7] <= 32'b00000000000000000000000000000000;
					memory[8] <= 32'b00000000000000000000000000000000;// BRANCH
					memory[9] <= 32'b00000000000000000000000000000000;
					memory[10] <= 32'b00000000000000000000000000000000;
					memory[11] <= 32'b00000000000000000000000000000000;
					memory[12] <= 32'b00000000000000000000000000000000;
					memory[13] <= 32'b00000000000000000000000000000000;
					memory[14] <= 32'b00000000000000000000000000000000;
					//memory[14] <= 32'b100011_00000_00000_0000000000000000;// LW
					/*memory[15] = 32'b00000000000000000000000000000000;
					memory[16] = 32'b00000000000000000000000000000000;
					memory[17] = 32'b00000000000000000000000000000000;
					memory[18] = 32'b00000000000000000000000000000000;
					memory[19] = 32'b00000000000000000000000000000000;///////////////////////////
					memory[20] = 32'b00000000000000000000000000000000;
					memory[21] = 32'b10001100000010110000000000000000;*/			
				end else begin
					for (j = 8'b0000_0100; j < 128; j = j + 8'b00000001) begin
						memory[j] <= 32'h0000_0000;
					end
					
					memory[0] <= 32'b00000000000000000000000000000010;
					memory[1] <= 32'b00000000000000000000000000000010;
					memory[2] <= 32'b00000000000000000000000000000010;
					memory[3] <= 32'b00000000000000000000000000000010;
					
				end
			end
    end

endmodule
