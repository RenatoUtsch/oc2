module Ram (
    input    [6:0]    addr,
    inout    [31:0]    data,
    input              wre,
	 input				  flag,	//memoria de dados/memoria de instrucoes
	 input 				  reset
);

    reg     [31:0]  memory    [0:127];
	 reg     [7:0] i;

    assign data[31:0] = wre ? memory[addr] : 32'hZZZZ_ZZZZ;

    always @(wre or addr or data or reset) begin
        if (!wre)
            memory[addr] = data[31:0];
				
			if(!reset) begin
				if(flag)begin			
				
					for (i = 0; i < 128; i = i + 1) begin
						memory[i] = 32'h0000_0000;
					end
					
					memory[0] = 32'b00000000000000000000000000000000;
					memory[1] = 32'b00000000000000000000000000000000;
					memory[2] = 32'b00000000000000000000000000000000;
					memory[3] = 32'b00001000000000000000000000001111;///////////////////////////
					memory[4] = 32'b00000000000000000000000000000000;
					memory[5] = 32'b00000000000000000000000000000000;
					memory[6] = 32'b00000000000000000000000000000000;
					memory[7] = 32'b00100000101001010000000000000101;///////////////////////////
					memory[8] = 32'b00000000000000000000000000000000;
					memory[9] = 32'b00000000000000000000000000000000;
					memory[10] = 32'b00000000000000000000000000000000;
					memory[11] = 32'b00010000100001011111111111110111;///////////////////////////
					memory[12] = 32'b00000000000000000000000000000000;
					memory[13] = 32'b00000000000000000000000000000000;
					memory[14] = 32'b00000000000000000000000000000000;
					memory[15] = 32'b00000000100001010011000000100000;///////////////////////////
					memory[16] = 32'b00000000000000000000000000000000;
					memory[17] = 32'b00000000000000000000000000000000;
					memory[18] = 32'b00000000000000000000000000000000;
					memory[19] = 32'b00100000000001110000000000001001;///////////////////////////
					memory[20] = 32'b00000000000000000000000000000000;
					memory[21] = 32'b00000000000000000000000000000000;
					
					
				end
			end
    end

endmodule
