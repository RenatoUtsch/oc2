module Execute_Y (
    input               clock,
    input               reset,
    // Issue
);

    Execute_Y0 e_Y0();
    Execute_Y1 e_Y1();
    Execute_Y2 e_Y2();
    Execute_Y3 e_Y3();

endmodule

module Execute_Y0 (

);



endmodule

module Execute_Y1 (

);



endmodule

module Execute_Y2 (

);



endmodule

module Execute_Y3 (

);



endmodule
